module encoder4x2(
  input [3:0]x,
  output reg [1:0]y);
  always@(*) begin
    case(x)
      4'b1000:assign y=2'b00;
      4'b0100:assign y=2'b01;
      4'b0010:assign y=2'b10;
      4'b0001:assign y=2'b11;
    endcase
  end
endmodule
